VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRF_2R1W
  CLASS BLOCK ;
  FOREIGN DFFRF_2R1W ;
  ORIGIN 0.000 0.000 ;
  SIZE 358.800 BY 176.800 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 2.000 88.360 ;
    END
  END CLK
  PIN DA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 174.800 3.130 176.800 ;
    END
  END DA[0]
  PIN DA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 174.800 58.790 176.800 ;
    END
  END DA[10]
  PIN DA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 174.800 64.770 176.800 ;
    END
  END DA[11]
  PIN DA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 174.800 70.290 176.800 ;
    END
  END DA[12]
  PIN DA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 174.800 75.810 176.800 ;
    END
  END DA[13]
  PIN DA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 174.800 81.330 176.800 ;
    END
  END DA[14]
  PIN DA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 174.800 86.850 176.800 ;
    END
  END DA[15]
  PIN DA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 174.800 92.830 176.800 ;
    END
  END DA[16]
  PIN DA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 174.800 98.350 176.800 ;
    END
  END DA[17]
  PIN DA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 174.800 103.870 176.800 ;
    END
  END DA[18]
  PIN DA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 174.800 109.390 176.800 ;
    END
  END DA[19]
  PIN DA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 174.800 8.650 176.800 ;
    END
  END DA[1]
  PIN DA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 174.800 114.910 176.800 ;
    END
  END DA[20]
  PIN DA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 174.800 120.430 176.800 ;
    END
  END DA[21]
  PIN DA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 174.800 126.410 176.800 ;
    END
  END DA[22]
  PIN DA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 174.800 131.930 176.800 ;
    END
  END DA[23]
  PIN DA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 174.800 137.450 176.800 ;
    END
  END DA[24]
  PIN DA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 174.800 142.970 176.800 ;
    END
  END DA[25]
  PIN DA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 174.800 148.490 176.800 ;
    END
  END DA[26]
  PIN DA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 174.800 154.470 176.800 ;
    END
  END DA[27]
  PIN DA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 174.800 159.990 176.800 ;
    END
  END DA[28]
  PIN DA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 174.800 165.510 176.800 ;
    END
  END DA[29]
  PIN DA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 174.800 14.170 176.800 ;
    END
  END DA[2]
  PIN DA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 174.800 171.030 176.800 ;
    END
  END DA[30]
  PIN DA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 174.800 176.550 176.800 ;
    END
  END DA[31]
  PIN DA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 174.800 19.690 176.800 ;
    END
  END DA[3]
  PIN DA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 174.800 25.210 176.800 ;
    END
  END DA[4]
  PIN DA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 174.800 30.730 176.800 ;
    END
  END DA[5]
  PIN DA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 174.800 36.710 176.800 ;
    END
  END DA[6]
  PIN DA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 174.800 42.230 176.800 ;
    END
  END DA[7]
  PIN DA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 174.800 47.750 176.800 ;
    END
  END DA[8]
  PIN DA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 174.800 53.270 176.800 ;
    END
  END DA[9]
  PIN DB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 174.800 182.530 176.800 ;
    END
  END DB[0]
  PIN DB[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 174.800 238.190 176.800 ;
    END
  END DB[10]
  PIN DB[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 174.800 244.170 176.800 ;
    END
  END DB[11]
  PIN DB[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 174.800 249.690 176.800 ;
    END
  END DB[12]
  PIN DB[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 174.800 255.210 176.800 ;
    END
  END DB[13]
  PIN DB[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 174.800 260.730 176.800 ;
    END
  END DB[14]
  PIN DB[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 174.800 266.250 176.800 ;
    END
  END DB[15]
  PIN DB[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 174.800 272.230 176.800 ;
    END
  END DB[16]
  PIN DB[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 174.800 277.750 176.800 ;
    END
  END DB[17]
  PIN DB[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 174.800 283.270 176.800 ;
    END
  END DB[18]
  PIN DB[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 174.800 288.790 176.800 ;
    END
  END DB[19]
  PIN DB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 174.800 188.050 176.800 ;
    END
  END DB[1]
  PIN DB[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 174.800 294.310 176.800 ;
    END
  END DB[20]
  PIN DB[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 174.800 299.830 176.800 ;
    END
  END DB[21]
  PIN DB[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 174.800 305.810 176.800 ;
    END
  END DB[22]
  PIN DB[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 174.800 311.330 176.800 ;
    END
  END DB[23]
  PIN DB[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 174.800 316.850 176.800 ;
    END
  END DB[24]
  PIN DB[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 174.800 322.370 176.800 ;
    END
  END DB[25]
  PIN DB[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 174.800 327.890 176.800 ;
    END
  END DB[26]
  PIN DB[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 174.800 333.870 176.800 ;
    END
  END DB[27]
  PIN DB[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 174.800 339.390 176.800 ;
    END
  END DB[28]
  PIN DB[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 174.800 344.910 176.800 ;
    END
  END DB[29]
  PIN DB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 174.800 193.570 176.800 ;
    END
  END DB[2]
  PIN DB[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 174.800 350.430 176.800 ;
    END
  END DB[30]
  PIN DB[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 174.800 355.950 176.800 ;
    END
  END DB[31]
  PIN DB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 174.800 199.090 176.800 ;
    END
  END DB[3]
  PIN DB[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 174.800 204.610 176.800 ;
    END
  END DB[4]
  PIN DB[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 174.800 210.130 176.800 ;
    END
  END DB[5]
  PIN DB[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 174.800 216.110 176.800 ;
    END
  END DB[6]
  PIN DB[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 174.800 221.630 176.800 ;
    END
  END DB[7]
  PIN DB[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 174.800 227.150 176.800 ;
    END
  END DB[8]
  PIN DB[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 174.800 232.670 176.800 ;
    END
  END DB[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.000 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.000 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 2.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 2.000 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 2.000 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 2.000 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 2.000 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 2.000 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 2.000 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 2.000 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 2.000 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.000 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 2.000 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 2.000 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 2.000 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 2.000 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 2.000 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 2.000 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 2.000 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 2.000 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 2.000 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 2.000 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.000 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 2.000 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 2.000 ;
    END
  END DW[31]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.000 ;
    END
  END DW[3]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.000 ;
    END
  END DW[4]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.000 ;
    END
  END DW[5]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.000 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.000 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.000 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 2.000 ;
    END
  END DW[9]
  PIN RA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 8.880 358.800 9.480 ;
    END
  END RA[0]
  PIN RA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 26.560 358.800 27.160 ;
    END
  END RA[1]
  PIN RA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 44.240 358.800 44.840 ;
    END
  END RA[2]
  PIN RA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 61.920 358.800 62.520 ;
    END
  END RA[3]
  PIN RA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 79.600 358.800 80.200 ;
    END
  END RA[4]
  PIN RB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 97.280 358.800 97.880 ;
    END
  END RB[0]
  PIN RB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 114.960 358.800 115.560 ;
    END
  END RB[1]
  PIN RB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 132.640 358.800 133.240 ;
    END
  END RB[2]
  PIN RB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 150.320 358.800 150.920 ;
    END
  END RB[3]
  PIN RB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.800 168.000 358.800 168.600 ;
    END
  END RB[4]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.000 12.880 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.000 38.040 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.000 63.200 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 2.000 138.680 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 2.000 163.840 ;
    END
  END RW[4]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 174.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 174.320 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 174.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 174.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 174.320 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.000 113.520 ;
    END
  END WE
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 356.040 174.165 ;
      LAYER met1 ;
        RECT 2.370 0.040 356.040 176.760 ;
      LAYER met2 ;
        RECT 2.400 174.520 2.570 176.790 ;
        RECT 3.410 174.520 8.090 176.790 ;
        RECT 8.930 174.520 13.610 176.790 ;
        RECT 14.450 174.520 19.130 176.790 ;
        RECT 19.970 174.520 24.650 176.790 ;
        RECT 25.490 174.520 30.170 176.790 ;
        RECT 31.010 174.520 36.150 176.790 ;
        RECT 36.990 174.520 41.670 176.790 ;
        RECT 42.510 174.520 47.190 176.790 ;
        RECT 48.030 174.520 52.710 176.790 ;
        RECT 53.550 174.520 58.230 176.790 ;
        RECT 59.070 174.520 64.210 176.790 ;
        RECT 65.050 174.520 69.730 176.790 ;
        RECT 70.570 174.520 75.250 176.790 ;
        RECT 76.090 174.520 80.770 176.790 ;
        RECT 81.610 174.520 86.290 176.790 ;
        RECT 87.130 174.520 92.270 176.790 ;
        RECT 93.110 174.520 97.790 176.790 ;
        RECT 98.630 174.520 103.310 176.790 ;
        RECT 104.150 174.520 108.830 176.790 ;
        RECT 109.670 174.520 114.350 176.790 ;
        RECT 115.190 174.520 119.870 176.790 ;
        RECT 120.710 174.520 125.850 176.790 ;
        RECT 126.690 174.520 131.370 176.790 ;
        RECT 132.210 174.520 136.890 176.790 ;
        RECT 137.730 174.520 142.410 176.790 ;
        RECT 143.250 174.520 147.930 176.790 ;
        RECT 148.770 174.520 153.910 176.790 ;
        RECT 154.750 174.520 159.430 176.790 ;
        RECT 160.270 174.520 164.950 176.790 ;
        RECT 165.790 174.520 170.470 176.790 ;
        RECT 171.310 174.520 175.990 176.790 ;
        RECT 176.830 174.520 181.970 176.790 ;
        RECT 182.810 174.520 187.490 176.790 ;
        RECT 188.330 174.520 193.010 176.790 ;
        RECT 193.850 174.520 198.530 176.790 ;
        RECT 199.370 174.520 204.050 176.790 ;
        RECT 204.890 174.520 209.570 176.790 ;
        RECT 210.410 174.520 215.550 176.790 ;
        RECT 216.390 174.520 221.070 176.790 ;
        RECT 221.910 174.520 226.590 176.790 ;
        RECT 227.430 174.520 232.110 176.790 ;
        RECT 232.950 174.520 237.630 176.790 ;
        RECT 238.470 174.520 243.610 176.790 ;
        RECT 244.450 174.520 249.130 176.790 ;
        RECT 249.970 174.520 254.650 176.790 ;
        RECT 255.490 174.520 260.170 176.790 ;
        RECT 261.010 174.520 265.690 176.790 ;
        RECT 266.530 174.520 271.670 176.790 ;
        RECT 272.510 174.520 277.190 176.790 ;
        RECT 278.030 174.520 282.710 176.790 ;
        RECT 283.550 174.520 288.230 176.790 ;
        RECT 289.070 174.520 293.750 176.790 ;
        RECT 294.590 174.520 299.270 176.790 ;
        RECT 300.110 174.520 305.250 176.790 ;
        RECT 306.090 174.520 310.770 176.790 ;
        RECT 311.610 174.520 316.290 176.790 ;
        RECT 317.130 174.520 321.810 176.790 ;
        RECT 322.650 174.520 327.330 176.790 ;
        RECT 328.170 174.520 333.310 176.790 ;
        RECT 334.150 174.520 338.830 176.790 ;
        RECT 339.670 174.520 344.350 176.790 ;
        RECT 345.190 174.520 349.870 176.790 ;
        RECT 350.710 174.520 355.390 176.790 ;
        RECT 2.400 2.280 355.940 174.520 ;
        RECT 2.400 0.010 5.330 2.280 ;
        RECT 6.170 0.010 16.370 2.280 ;
        RECT 17.210 0.010 27.410 2.280 ;
        RECT 28.250 0.010 38.910 2.280 ;
        RECT 39.750 0.010 49.950 2.280 ;
        RECT 50.790 0.010 60.990 2.280 ;
        RECT 61.830 0.010 72.490 2.280 ;
        RECT 73.330 0.010 83.530 2.280 ;
        RECT 84.370 0.010 95.030 2.280 ;
        RECT 95.870 0.010 106.070 2.280 ;
        RECT 106.910 0.010 117.110 2.280 ;
        RECT 117.950 0.010 128.610 2.280 ;
        RECT 129.450 0.010 139.650 2.280 ;
        RECT 140.490 0.010 150.690 2.280 ;
        RECT 151.530 0.010 162.190 2.280 ;
        RECT 163.030 0.010 173.230 2.280 ;
        RECT 174.070 0.010 184.730 2.280 ;
        RECT 185.570 0.010 195.770 2.280 ;
        RECT 196.610 0.010 206.810 2.280 ;
        RECT 207.650 0.010 218.310 2.280 ;
        RECT 219.150 0.010 229.350 2.280 ;
        RECT 230.190 0.010 240.390 2.280 ;
        RECT 241.230 0.010 251.890 2.280 ;
        RECT 252.730 0.010 262.930 2.280 ;
        RECT 263.770 0.010 274.430 2.280 ;
        RECT 275.270 0.010 285.470 2.280 ;
        RECT 286.310 0.010 296.510 2.280 ;
        RECT 297.350 0.010 308.010 2.280 ;
        RECT 308.850 0.010 319.050 2.280 ;
        RECT 319.890 0.010 330.090 2.280 ;
        RECT 330.930 0.010 341.590 2.280 ;
        RECT 342.430 0.010 352.630 2.280 ;
        RECT 353.470 0.010 355.940 2.280 ;
      LAYER met3 ;
        RECT 2.000 169.000 356.800 176.625 ;
        RECT 2.000 167.600 356.400 169.000 ;
        RECT 2.000 164.240 356.800 167.600 ;
        RECT 2.400 162.840 356.800 164.240 ;
        RECT 2.000 151.320 356.800 162.840 ;
        RECT 2.000 149.920 356.400 151.320 ;
        RECT 2.000 139.080 356.800 149.920 ;
        RECT 2.400 137.680 356.800 139.080 ;
        RECT 2.000 133.640 356.800 137.680 ;
        RECT 2.000 132.240 356.400 133.640 ;
        RECT 2.000 115.960 356.800 132.240 ;
        RECT 2.000 114.560 356.400 115.960 ;
        RECT 2.000 113.920 356.800 114.560 ;
        RECT 2.400 112.520 356.800 113.920 ;
        RECT 2.000 98.280 356.800 112.520 ;
        RECT 2.000 96.880 356.400 98.280 ;
        RECT 2.000 88.760 356.800 96.880 ;
        RECT 2.400 87.360 356.800 88.760 ;
        RECT 2.000 80.600 356.800 87.360 ;
        RECT 2.000 79.200 356.400 80.600 ;
        RECT 2.000 63.600 356.800 79.200 ;
        RECT 2.400 62.920 356.800 63.600 ;
        RECT 2.400 62.200 356.400 62.920 ;
        RECT 2.000 61.520 356.400 62.200 ;
        RECT 2.000 45.240 356.800 61.520 ;
        RECT 2.000 43.840 356.400 45.240 ;
        RECT 2.000 38.440 356.800 43.840 ;
        RECT 2.400 37.040 356.800 38.440 ;
        RECT 2.000 27.560 356.800 37.040 ;
        RECT 2.000 26.160 356.400 27.560 ;
        RECT 2.000 13.280 356.800 26.160 ;
        RECT 2.400 11.880 356.800 13.280 ;
        RECT 2.000 9.880 356.800 11.880 ;
        RECT 2.000 8.480 356.400 9.880 ;
        RECT 2.000 0.175 356.800 8.480 ;
      LAYER met4 ;
        RECT 93.215 174.720 344.705 176.625 ;
        RECT 93.215 19.895 94.680 174.720 ;
        RECT 97.080 19.895 171.480 174.720 ;
        RECT 173.880 19.895 248.280 174.720 ;
        RECT 250.680 19.895 325.080 174.720 ;
        RECT 327.480 19.895 344.705 174.720 ;
  END
END DFFRF_2R1W
END LIBRARY

