VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32
  CLASS BLOCK ;
  FOREIGN RAM32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 399.280 BY 100.640 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 55.120 399.280 55.720 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 64.640 399.280 65.240 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 74.840 399.280 75.440 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 85.040 399.280 85.640 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 95.240 399.280 95.840 ;
    END
  END A0[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.000 50.960 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 98.640 6.350 100.640 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 98.640 131.010 100.640 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 98.640 143.430 100.640 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 98.640 155.850 100.640 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 98.640 168.270 100.640 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 98.640 180.690 100.640 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 98.640 193.110 100.640 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 98.640 205.990 100.640 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 98.640 218.410 100.640 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 98.640 230.830 100.640 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 98.640 243.250 100.640 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 98.640 18.770 100.640 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 98.640 255.670 100.640 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 98.640 268.090 100.640 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 98.640 280.510 100.640 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 98.640 292.930 100.640 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 98.640 305.810 100.640 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 98.640 318.230 100.640 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 98.640 330.650 100.640 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 98.640 343.070 100.640 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 98.640 355.490 100.640 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 98.640 367.910 100.640 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 98.640 31.190 100.640 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 98.640 380.330 100.640 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 98.640 392.750 100.640 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 98.640 43.610 100.640 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 98.640 56.030 100.640 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 98.640 68.450 100.640 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 98.640 80.870 100.640 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 98.640 93.290 100.640 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 98.640 106.170 100.640 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 98.640 118.590 100.640 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 4.800 399.280 5.400 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 98.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 98.160 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 14.320 399.280 14.920 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 24.520 399.280 25.120 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 34.720 399.280 35.320 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.280 44.920 399.280 45.520 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 396.520 98.005 ;
      LAYER met1 ;
        RECT 2.760 0.380 396.520 100.600 ;
      LAYER met2 ;
        RECT 4.700 98.360 5.790 100.630 ;
        RECT 6.630 98.360 18.210 100.630 ;
        RECT 19.050 98.360 30.630 100.630 ;
        RECT 31.470 98.360 43.050 100.630 ;
        RECT 43.890 98.360 55.470 100.630 ;
        RECT 56.310 98.360 67.890 100.630 ;
        RECT 68.730 98.360 80.310 100.630 ;
        RECT 81.150 98.360 92.730 100.630 ;
        RECT 93.570 98.360 105.610 100.630 ;
        RECT 106.450 98.360 118.030 100.630 ;
        RECT 118.870 98.360 130.450 100.630 ;
        RECT 131.290 98.360 142.870 100.630 ;
        RECT 143.710 98.360 155.290 100.630 ;
        RECT 156.130 98.360 167.710 100.630 ;
        RECT 168.550 98.360 180.130 100.630 ;
        RECT 180.970 98.360 192.550 100.630 ;
        RECT 193.390 98.360 205.430 100.630 ;
        RECT 206.270 98.360 217.850 100.630 ;
        RECT 218.690 98.360 230.270 100.630 ;
        RECT 231.110 98.360 242.690 100.630 ;
        RECT 243.530 98.360 255.110 100.630 ;
        RECT 255.950 98.360 267.530 100.630 ;
        RECT 268.370 98.360 279.950 100.630 ;
        RECT 280.790 98.360 292.370 100.630 ;
        RECT 293.210 98.360 305.250 100.630 ;
        RECT 306.090 98.360 317.670 100.630 ;
        RECT 318.510 98.360 330.090 100.630 ;
        RECT 330.930 98.360 342.510 100.630 ;
        RECT 343.350 98.360 354.930 100.630 ;
        RECT 355.770 98.360 367.350 100.630 ;
        RECT 368.190 98.360 379.770 100.630 ;
        RECT 380.610 98.360 392.190 100.630 ;
        RECT 393.030 98.360 396.430 100.630 ;
        RECT 4.700 2.280 396.430 98.360 ;
        RECT 4.700 0.155 5.790 2.280 ;
        RECT 6.630 0.155 18.210 2.280 ;
        RECT 19.050 0.155 30.630 2.280 ;
        RECT 31.470 0.155 43.050 2.280 ;
        RECT 43.890 0.155 55.470 2.280 ;
        RECT 56.310 0.155 67.890 2.280 ;
        RECT 68.730 0.155 80.310 2.280 ;
        RECT 81.150 0.155 92.730 2.280 ;
        RECT 93.570 0.155 105.610 2.280 ;
        RECT 106.450 0.155 118.030 2.280 ;
        RECT 118.870 0.155 130.450 2.280 ;
        RECT 131.290 0.155 142.870 2.280 ;
        RECT 143.710 0.155 155.290 2.280 ;
        RECT 156.130 0.155 167.710 2.280 ;
        RECT 168.550 0.155 180.130 2.280 ;
        RECT 180.970 0.155 192.550 2.280 ;
        RECT 193.390 0.155 205.430 2.280 ;
        RECT 206.270 0.155 217.850 2.280 ;
        RECT 218.690 0.155 230.270 2.280 ;
        RECT 231.110 0.155 242.690 2.280 ;
        RECT 243.530 0.155 255.110 2.280 ;
        RECT 255.950 0.155 267.530 2.280 ;
        RECT 268.370 0.155 279.950 2.280 ;
        RECT 280.790 0.155 292.370 2.280 ;
        RECT 293.210 0.155 305.250 2.280 ;
        RECT 306.090 0.155 317.670 2.280 ;
        RECT 318.510 0.155 330.090 2.280 ;
        RECT 330.930 0.155 342.510 2.280 ;
        RECT 343.350 0.155 354.930 2.280 ;
        RECT 355.770 0.155 367.350 2.280 ;
        RECT 368.190 0.155 379.770 2.280 ;
        RECT 380.610 0.155 392.190 2.280 ;
        RECT 393.030 0.155 396.430 2.280 ;
      LAYER met3 ;
        RECT 2.000 96.240 397.280 99.785 ;
        RECT 2.000 94.840 396.880 96.240 ;
        RECT 2.000 86.040 397.280 94.840 ;
        RECT 2.000 84.640 396.880 86.040 ;
        RECT 2.000 75.840 397.280 84.640 ;
        RECT 2.000 74.440 396.880 75.840 ;
        RECT 2.000 65.640 397.280 74.440 ;
        RECT 2.000 64.240 396.880 65.640 ;
        RECT 2.000 56.120 397.280 64.240 ;
        RECT 2.000 54.720 396.880 56.120 ;
        RECT 2.000 51.360 397.280 54.720 ;
        RECT 2.400 49.960 397.280 51.360 ;
        RECT 2.000 45.920 397.280 49.960 ;
        RECT 2.000 44.520 396.880 45.920 ;
        RECT 2.000 35.720 397.280 44.520 ;
        RECT 2.000 34.320 396.880 35.720 ;
        RECT 2.000 25.520 397.280 34.320 ;
        RECT 2.000 24.120 396.880 25.520 ;
        RECT 2.000 15.320 397.280 24.120 ;
        RECT 2.000 13.920 396.880 15.320 ;
        RECT 2.000 5.800 397.280 13.920 ;
        RECT 2.000 4.400 396.880 5.800 ;
        RECT 2.000 0.175 397.280 4.400 ;
      LAYER met4 ;
        RECT 111.615 28.735 111.945 31.785 ;
  END
END RAM32
END LIBRARY

